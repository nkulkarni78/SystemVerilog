interface d_intf();
  logic reset;
  logic [3:0]d;
  logic [3:0]q;
  logic clock;
endinterface
