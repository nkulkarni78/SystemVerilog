interface d_intf();
  logic tb_reset;
  logic [3:0]tb_d;
  logic [3:0]tb_q;
  logic clock;
endinterface
